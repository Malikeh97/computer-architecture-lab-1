module IF_Stage(
	input clk,
	input rst,
	input Br_tacken,
	input[31:0] Br_Addr,
	output[31:0] PC,
	output[31:0] Instruction
);

reg[31:0] pc = 32'b0;
reg[31:0] ROM[127:0];

initial begin
	ROM[0]  <= 32'b10000000000000010000011000001010;
	ROM[1]  <= 32'b00000100000000010001000000000000;
	ROM[2]  <= 32'b00001100000000010001100000000000;
	ROM[3]  <= 32'b00010100010000110010000000000000;
	ROM[4]  <= 32'b10000100011001010001101000110100;
	ROM[5]  <= 32'b00011000011001000010100000000000;
	ROM[6]  <= 32'b00011100101000000011000000000000;
	ROM[7]  <= 32'b00011100100000000101100000000000;
	ROM[8]  <= 32'b00001100101001010010100000000000;
	ROM[9]  <= 32'b10000000000000010000010000000000;
	ROM[10] <= 32'b10010100001000100000000000000000;
	ROM[11] <= 32'b10010000001001010000000000000000;
	ROM[12] <= 32'b10100000101000000000000000000001;
	ROM[13] <= 32'b00100000101000010011100000000000;
	ROM[14] <= 32'b00100000101000010000000000000000;
	ROM[15] <= 32'b00100100011010110011100000000000;
	ROM[16] <= 32'b00101000011010110100000000000000;
	ROM[17] <= 32'b00101100011001000100100000000000;
	ROM[18] <= 32'b00110000011001000101000000000000;
	ROM[19] <= 32'b10010100001000110000000000000100;
	ROM[20] <= 32'b10010100001001000000000000001000;
	ROM[21] <= 32'b10010100001001010000000000001100;
	ROM[22] <= 32'b10010100001001100000000000010000;
	ROM[23] <= 32'b10010000001010110000000000000100;
	ROM[24] <= 32'b10010100001001110000000000010100;
	ROM[25] <= 32'b10010100001010000000000000011000;
	ROM[26] <= 32'b10010100001010010000000000011100;
	ROM[27] <= 32'b10010100001010100000000000100000;
	ROM[28] <= 32'b10010100001010110000000000100100;
	ROM[29] <= 32'b10000000000000010000000000000011;
	ROM[30] <= 32'b10000000000001000000010000000000;
	ROM[31] <= 32'b10000000000000100000000000000000;
	ROM[32] <= 32'b10000000000000110000000000000001;
	ROM[33] <= 32'b10000000000010010000000000000010;
	ROM[34] <= 32'b00101000011010010100000000000000;
	ROM[35] <= 32'b00000100100010000100000000000000;
	ROM[36] <= 32'b10010001000001010000000000000000;
	ROM[37] <= 32'b10010001000001101111111111111100;
	ROM[38] <= 32'b00001100101001100100100000000000;
	ROM[39] <= 32'b10000000000010101000000000000000;
	ROM[40] <= 32'b10000000000010110000000000010000;
	ROM[41] <= 32'b00101001010010110101000000000000;
	ROM[42] <= 32'b00010101001010100100100000000000;
	ROM[43] <= 32'b10100001001000000000000000000010;
	ROM[44] <= 32'b10010101000001011111111111111100;
	ROM[45] <= 32'b10010101000001100000000000000000;
	ROM[46] <= 32'b10000000011000110000000000000001;
	ROM[47] <= 32'b10100100001000111111111111110001;
	ROM[48] <= 32'b10000000010000100000000000000001;
	ROM[49] <= 32'b10100100001000101111111111101110;
	ROM[50] <= 32'b10000000000000010000010000000000;
	ROM[51] <= 32'b10010000001000100000000000000000;
	ROM[52] <= 32'b10010000001000110000000000000100;
	ROM[53] <= 32'b10010000001001000000000000001000;
	ROM[54] <= 32'b10010000001001000000001000001000;
	ROM[55] <= 32'b10010000001001000000010000001000;
	ROM[56] <= 32'b10010000001001010000000000001100;
	ROM[57] <= 32'b10010000001001100000000000010000;
	ROM[58] <= 32'b10010000001001110000000000010100;
	ROM[59] <= 32'b10010000001010000000000000011000;
	ROM[60] <= 32'b10010000001010010000000000011100;
	ROM[61] <= 32'b10010000001010100000000000100000;
	ROM[62] <= 32'b10010000001010110000000000100100;
	ROM[63] <= 32'b10101000000000001111111111111111;
end

always  @(posedge clk, posedge rst)begin
	if(rst) pc <= 32'b0;
	else pc <= Br_tacken ? Br_Addr: pc + 32'd4;
end

assign PC = pc;
assign Instruction = ROM[PC[31:2]];

endmodule
